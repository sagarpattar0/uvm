module simpand(input wire clk,
                input wire en,
                input wire a,
                input wire b,
                 output reg y);




