`include "uvm_macros.svh"
import uvm_pkg::*;

interface simpleand_inf;
  logic a;
  logic b;
  logic y;
  logic clk;
  logic en;
endinterface: simpleand_inf
